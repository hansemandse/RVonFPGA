-- ***********************************************************************
--              |
-- Title        : Implementation and Optimization of a RISC-V Processor on
--              : a FPGA
--              |
-- Developers   : Hans Jakob Damsgaard, Technical University of Denmark
--              : s163915@student.dtu.dk or hansjakobdamsgaard@gmail.com
--              |
-- Purpose      : This file is a part of a full system implemented as part
--              : of a bachelor's thesis at DTU. The thesis is written in
--              : cooperation with the Institute of Mathematics and
--              : Computer Science.
--              : This entity is a generated ROM containing the bootloader
--              : from the compiler.
--              |
-- Revision     : 1.0   (last updated June 28, 2019)
--              |
-- Available at : https://github.com/hansemandse/RVonFPGA
--              |
-- ***********************************************************************

library IEEE;
use IEEE.std_logic_1164.all;

library work;
use work.includes.all;

entity rom_gen is
    port (
        clk, reset : in std_logic;
        -- Memory interface
        Addr : in std_logic_vector(11 downto 0);
        ReadData : out std_logic_vector(DATA_WIDTH-1 downto 0)
    );
end rom_gen;

architecture rtl of rom_gen is
begin
    process (all)
    begin
        if (rising_edge(clk)) then
            if (reset = '1') then
                ReadData <= (others => '0');
            else
                case (Addr) is
					when x"000" => ReadData <= x"0b8000ef00000513";
					when x"008" => ReadData <= x"0010011b0a0000ef";
					when x"010" => ReadData <= x"00f1011303011113";
					when x"018" => ReadData <= x"0000119700c11113";
					when x"020" => ReadData <= x"0dc000ef6e418193";
					when x"028" => ReadData <= x"03c595930010059b";
					when x"030" => ReadData <= x"0005006700b56533";
					when x"038" => ReadData <= x"03f51513fff00513";
					when x"040" => ReadData <= x"0005050300350513";
					when x"048" => ReadData <= x"000080670ff57513";
					when x"050" => ReadData <= x"03f51513fff00513";
					when x"058" => ReadData <= x"0005050300250513";
					when x"060" => ReadData <= x"000080670ff57513";
					when x"068" => ReadData <= x"03f51513fff00513";
					when x"070" => ReadData <= x"0007878300350793";
					when x"078" => ReadData <= x"000794630ff7f793";
					when x"080" => ReadData <= x"001505130000006f";
					when x"088" => ReadData <= x"0ff5751300050503";
					when x"090" => ReadData <= x"fff0079300008067";
					when x"098" => ReadData <= x"0017879303f79793";
					when x"0a0" => ReadData <= x"0000806700a78023";
					when x"0a8" => ReadData <= x"03f79793fff00793";
					when x"0b0" => ReadData <= x"00a7802300478793";
					when x"0b8" => ReadData <= x"fff0079300008067";
					when x"0c0" => ReadData <= x"0057879303f79793";
					when x"0c8" => ReadData <= x"0000806700a78023";
					when x"0d0" => ReadData <= x"03f51513fff00513";
					when x"0d8" => ReadData <= x"0005050300450513";
					when x"0e0" => ReadData <= x"000080670ff57513";
					when x"0e8" => ReadData <= x"03f51513fff00513";
					when x"0f0" => ReadData <= x"0005050300550513";
					when x"0f8" => ReadData <= x"000080670ff57513";
					when x"100" => ReadData <= x"03f89893fff00893";
					when x"108" => ReadData <= x"00188e93f7010113";
					when x"110" => ReadData <= x"0ff37313000e8303";
					when x"118" => ReadData <= x"07213c2308913023";
					when x"120" => ReadData <= x"00001937fcf30f9b";
					when x"128" => ReadData <= x"fc930f1b000014b7";
					when x"130" => ReadData <= x"f00938030fffff93";
					when x"138" => ReadData <= x"0fff7f13f084be03";
					when x"140" => ReadData <= x"7f000793002f9293";
					when x"148" => ReadData <= x"0731382308813423";
					when x"150" => ReadData <= x"0751302307413423";
					when x"158" => ReadData <= x"0571382305613c23";
					when x"160" => ReadData <= x"0003039300100413";
					when x"168" => ReadData <= x"000f051300030593";
					when x"170" => ReadData <= x"0038879300f282b3";
					when x"178" => ReadData <= x"00078783000e8703";
					when x"180" => ReadData <= x"0ff7f7930ff77713";
					when x"188" => ReadData <= x"0007946305300693";
					when x"190" => ReadData <= x"fed71ce30000006f";
					when x"198" => ReadData <= x"0007878300388793";
					when x"1a0" => ReadData <= x"000794630ff7f793";
					when x"1a8" => ReadData <= x"fd03079b0000006f";
					when x"1b0" => ReadData <= x"009007130ff7f793";
					when x"1b8" => ReadData <= x"0390079362f76063";
					when x"1c0" => ReadData <= x"0077e663000f0713";
					when x"1c8" => ReadData <= x"0ff77713fd03871b";
					when x"1d0" => ReadData <= x"00e1002300388793";
					when x"1d8" => ReadData <= x"0ff7f79300078783";
					when x"1e0" => ReadData <= x"0000006f00079463";
					when x"1e8" => ReadData <= x"03900693000e8783";
					when x"1f0" => ReadData <= x"3ef6e8630ff7f793";
					when x"1f8" => ReadData <= x"0ff7f793fd07879b";
					when x"200" => ReadData <= x"0137e9b300471993";
					when x"208" => ReadData <= x"00f100a30019999b";
					when x"210" => ReadData <= x"080988630ff9f993";
					when x"218" => ReadData <= x"020a1a93fff98a1b";
					when x"220" => ReadData <= x"0001071300110693";
					when x"228" => ReadData <= x"fd058b9b020ada93";
					when x"230" => ReadData <= x"01568ab300388793";
					when x"238" => ReadData <= x"0007069300078783";
					when x"240" => ReadData <= x"03900b130ff7f793";
					when x"248" => ReadData <= x"000794630ffbfb93";
					when x"250" => ReadData <= x"000506130000006f";
					when x"258" => ReadData <= x"000b861300bb6463";
					when x"260" => ReadData <= x"0016869300c68023";
					when x"268" => ReadData <= x"001a5a1bff5692e3";
					when x"270" => ReadData <= x"00270693001a1a13";
					when x"278" => ReadData <= x"0080006f00da0a33";
					when x"280" => ReadData <= x"0007460300268693";
					when x"288" => ReadData <= x"0046161b00174783";
					when x"290" => ReadData <= x"00c7e7b300f7f793";
					when x"298" => ReadData <= x"0006871300f70023";
					when x"2a0" => ReadData <= x"0019d993ff4690e3";
					when x"2a8" => ReadData <= x"fff6071b0009861b";
					when x"2b0" => ReadData <= x"50d058630007069b";
					when x"2b8" => ReadData <= x"00c00a13ffe6079b";
					when x"2c0" => ReadData <= x"0037571b50fa7663";
					when x"2c8" => ReadData <= x"0001378300100a13";
					when x"2d0" => ReadData <= x"00813a0313470263";
					when x"2d8" => ReadData <= x"00200b130107fab3";
					when x"2e0" => ReadData <= x"010a7a330147c7b3";
					when x"2e8" => ReadData <= x"01c7f7b3014a8a33";
					when x"2f0" => ReadData <= x"1167006300fa47b3";
					when x"2f8" => ReadData <= x"0107fb3301013a03";
					when x"300" => ReadData <= x"00fa47b300300a93";
					when x"308" => ReadData <= x"016a0a33010a7a33";
					when x"310" => ReadData <= x"00fa47b301c7f7b3";
					when x"318" => ReadData <= x"01813a030d570e63";
					when x"320" => ReadData <= x"00400b130107fab3";
					when x"328" => ReadData <= x"010a7a3300fa47b3";
					when x"330" => ReadData <= x"01c7f7b3014a8a33";
					when x"338" => ReadData <= x"0b670c6300fa47b3";
					when x"340" => ReadData <= x"0107fab302013a03";
					when x"348" => ReadData <= x"0147c7b300500b13";
					when x"350" => ReadData <= x"014a8a33010a7a33";
					when x"358" => ReadData <= x"00fa47b301c7f7b3";
					when x"360" => ReadData <= x"02813a0309670a63";
					when x"368" => ReadData <= x"00600b130107fab3";
					when x"370" => ReadData <= x"010a7a330147c7b3";
					when x"378" => ReadData <= x"01c7f7b3014a8a33";
					when x"380" => ReadData <= x"0767086300fa47b3";
					when x"388" => ReadData <= x"0107fab303013a03";
					when x"390" => ReadData <= x"0147c7b300700b13";
					when x"398" => ReadData <= x"014a8a33010a7a33";
					when x"3a0" => ReadData <= x"00fa47b301c7f7b3";
					when x"3a8" => ReadData <= x"03813a0305670663";
					when x"3b0" => ReadData <= x"00800b130107fab3";
					when x"3b8" => ReadData <= x"010a7a330147c7b3";
					when x"3c0" => ReadData <= x"01c7f7b3014a8a33";
					when x"3c8" => ReadData <= x"0367046300fa47b3";
					when x"3d0" => ReadData <= x"f0093a8304013703";
					when x"3d8" => ReadData <= x"00e7ca33f084bb03";
					when x"3e0" => ReadData <= x"015777330157f7b3";
					when x"3e8" => ReadData <= x"016a77b300e78733";
					when x"3f0" => ReadData <= x"0087d71300f747b3";
					when x"3f8" => ReadData <= x"0107da1300f7073b";
					when x"400" => ReadData <= x"0147073b0137073b";
					when x"408" => ReadData <= x"0147073b0187da13";
					when x"410" => ReadData <= x"0147073b0207da13";
					when x"418" => ReadData <= x"0147073b0287da13";
					when x"420" => ReadData <= x"0147073b0307da13";
					when x"428" => ReadData <= x"00f707bb0387d793";
					when x"430" => ReadData <= x"0ff7f793ff86fa13";
					when x"438" => ReadData <= x"17468263000a071b";
					when x"440" => ReadData <= x"00ea0a3305010a13";
					when x"448" => ReadData <= x"00170a1bfb0a4a83";
					when x"450" => ReadData <= x"0ff7f79300fa87bb";
					when x"458" => ReadData <= x"05010a9314da5463";
					when x"460" => ReadData <= x"fb0a4a83014a8a33";
					when x"468" => ReadData <= x"00fa87bb00270a1b";
					when x"470" => ReadData <= x"12da56630ff7f793";
					when x"478" => ReadData <= x"014a8a3305010a93";
					when x"480" => ReadData <= x"00370a1bfb0a4a83";
					when x"488" => ReadData <= x"0ff7f79300fa87bb";
					when x"490" => ReadData <= x"05010a9310da5863";
					when x"498" => ReadData <= x"fb0a4a83014a8a33";
					when x"4a0" => ReadData <= x"00fa87bb00470a1b";
					when x"4a8" => ReadData <= x"0eda5a630ff7f793";
					when x"4b0" => ReadData <= x"014a8a3305010a93";
					when x"4b8" => ReadData <= x"00570a1bfb0a4a83";
					when x"4c0" => ReadData <= x"0ff7f79300fa87bb";
					when x"4c8" => ReadData <= x"05010a930cda5c63";
					when x"4d0" => ReadData <= x"fb0a4a83014a8a33";
					when x"4d8" => ReadData <= x"00fa87bb00670a1b";
					when x"4e0" => ReadData <= x"0ada5e630ff7f793";
					when x"4e8" => ReadData <= x"014a8a3305010a93";
					when x"4f0" => ReadData <= x"00770a1bfb0a4a83";
					when x"4f8" => ReadData <= x"0ff7f79300fa87bb";
					when x"500" => ReadData <= x"05010a930ada5063";
					when x"508" => ReadData <= x"fb0a4a83014a8a33";
					when x"510" => ReadData <= x"00fa87bb00870a1b";
					when x"518" => ReadData <= x"08da52630ff7f793";
					when x"520" => ReadData <= x"014a8a3305010a93";
					when x"528" => ReadData <= x"00970a1bfb0a4a83";
					when x"530" => ReadData <= x"0ff7f79300fa87bb";
					when x"538" => ReadData <= x"05010a9306da5463";
					when x"540" => ReadData <= x"fb0a4a83014a8a33";
					when x"548" => ReadData <= x"00fa87bb00a70a1b";
					when x"550" => ReadData <= x"04da56630ff7f793";
					when x"558" => ReadData <= x"014a8a3305010a93";
					when x"560" => ReadData <= x"00b70a1bfb0a4a83";
					when x"568" => ReadData <= x"0ff7f79300fa87bb";
					when x"570" => ReadData <= x"05010a9302da5863";
					when x"578" => ReadData <= x"fb0a4a03014a8a33";
					when x"580" => ReadData <= x"00fa07bb00c7071b";
					when x"588" => ReadData <= x"00d75a630ff7f793";
					when x"590" => ReadData <= x"fb07470300ea8733";
					when x"598" => ReadData <= x"0ff7f79300f707bb";
					when x"5a0" => ReadData <= x"00c7063305010713";
					when x"5a8" => ReadData <= x"fff74713fb064703";
					when x"5b0" => ReadData <= x"22f716630ff77713";
					when x"5b8" => ReadData <= x"03f7e06300800793";
					when x"5c0" => ReadData <= x"000780670002a783";
					when x"5c8" => ReadData <= x"0011468300014703";
					when x"5d0" => ReadData <= x"00d70733ffe4079b";
					when x"5d8" => ReadData <= x"0014041b20f71863";
					when x"5e0" => ReadData <= x"fc97879bb95ff06f";
					when x"5e8" => ReadData <= x"c15ff06f0ff7f793";
					when x"5f0" => ReadData <= x"0011470300014503";
					when x"5f8" => ReadData <= x"0021478300314683";
					when x"600" => ReadData <= x"0107171b0185151b";
					when x"608" => ReadData <= x"00d5653300e56533";
					when x"610" => ReadData <= x"00f565330087979b";
					when x"618" => ReadData <= x"088134030005051b";
					when x"620" => ReadData <= x"0781390308013483";
					when x"628" => ReadData <= x"06813a0307013983";
					when x"630" => ReadData <= x"05813b0306013a83";
					when x"638" => ReadData <= x"0901011305013b83";
					when x"640" => ReadData <= x"0001450300008067";
					when x"648" => ReadData <= x"0021470300114783";
					when x"650" => ReadData <= x"0087979b0105151b";
					when x"658" => ReadData <= x"00e5653300f56533";
					when x"660" => ReadData <= x"00015783fbdff06f";
					when x"668" => ReadData <= x"0087951b0087d71b";
					when x"670" => ReadData <= x"0305151300e56533";
					when x"678" => ReadData <= x"fa1ff06f03055513";
					when x"680" => ReadData <= x"0011470300014603";
					when x"688" => ReadData <= x"0021478300314a03";
					when x"690" => ReadData <= x"0107171b0186161b";
					when x"698" => ReadData <= x"0087979b00e66633";
					when x"6a0" => ReadData <= x"00f6663301466633";
					when x"6a8" => ReadData <= x"0006061b00400793";
					when x"6b0" => ReadData <= x"ffa9871bf2d7d6e3";
					when x"6b8" => ReadData <= x"0207571302071713";
					when x"6c0" => ReadData <= x"0011069300010793";
					when x"6c8" => ReadData <= x"00d7073300100a13";
					when x"6d0" => ReadData <= x"03ca1a1340f60633";
					when x"6d8" => ReadData <= x"0047c98300f606b3";
					when x"6e0" => ReadData <= x"013680230146e6b3";
					when x"6e8" => ReadData <= x"fee796e300178793";
					when x"6f0" => ReadData <= x"a81ff06f0014041b";
					when x"6f8" => ReadData <= x"0011478300014603";
					when x"700" => ReadData <= x"0106161b00214703";
					when x"708" => ReadData <= x"00f666330087979b";
					when x"710" => ReadData <= x"00e6663300300793";
					when x"718" => ReadData <= x"ffb9899becd7d2e3";
					when x"720" => ReadData <= x"0209d99302099993";
					when x"728" => ReadData <= x"0011071300010793";
					when x"730" => ReadData <= x"00e989b300100a13";
					when x"738" => ReadData <= x"03ca1a1340f60633";
					when x"740" => ReadData <= x"0037c68300f60733";
					when x"748" => ReadData <= x"00d7002301476733";
					when x"750" => ReadData <= x"ff3796e300178793";
					when x"758" => ReadData <= x"a19ff06f0014041b";
					when x"760" => ReadData <= x"0020071300015783";
					when x"768" => ReadData <= x"0087961b0087da1b";
					when x"770" => ReadData <= x"0306161301466633";
					when x"778" => ReadData <= x"e6d750e303065613";
					when x"780" => ReadData <= x"02099993ffc9899b";
					when x"788" => ReadData <= x"000107930209d993";
					when x"790" => ReadData <= x"00100a1300110713";
					when x"798" => ReadData <= x"40f6063300e989b3";
					when x"7a0" => ReadData <= x"00f6073303ca1a13";
					when x"7a8" => ReadData <= x"014767330027c683";
					when x"7b0" => ReadData <= x"0017879300d70023";
					when x"7b8" => ReadData <= x"0014041bff3796e3";
					when x"7c0" => ReadData <= x"000987939b5ff06f";
					when x"7c8" => ReadData <= x"00098793dd9ff06f";
					when x"7d0" => ReadData <= x"c6dff06f00000713";
					when x"7d8" => ReadData <= x"e41ff06ffff00513";
					when x"7e0" => ReadData <= x"e39ff06f00200513";
					when x"7e8" => ReadData <= x"e31ff06f00300513";
					when x"7f0" => ReadData <= x"000006f800000760";
					when x"7f8" => ReadData <= x"000005dc00000680";
					when x"800" => ReadData <= x"000005dc000005c8";
					when x"808" => ReadData <= x"0000064400000664";
					when x"810" => ReadData <= x"00000000000005f0";
					when x"818" => ReadData <= x"0000000000000000";
					when x"820" => ReadData <= x"0000000000000000";
					when x"828" => ReadData <= x"0000000000000000";
					when x"830" => ReadData <= x"0000000000000000";
					when x"838" => ReadData <= x"0000000000000000";
					when x"840" => ReadData <= x"0000000000000000";
					when x"848" => ReadData <= x"0000000000000000";
					when x"850" => ReadData <= x"0000000000000000";
					when x"858" => ReadData <= x"0000000000000000";
					when x"860" => ReadData <= x"0000000000000000";
					when x"868" => ReadData <= x"0000000000000000";
					when x"870" => ReadData <= x"0000000000000000";
					when x"878" => ReadData <= x"0000000000000000";
					when x"880" => ReadData <= x"0000000000000000";
					when x"888" => ReadData <= x"0000000000000000";
					when x"890" => ReadData <= x"0000000000000000";
					when x"898" => ReadData <= x"0000000000000000";
					when x"8a0" => ReadData <= x"0000000000000000";
					when x"8a8" => ReadData <= x"0000000000000000";
					when x"8b0" => ReadData <= x"0000000000000000";
					when x"8b8" => ReadData <= x"0000000000000000";
					when x"8c0" => ReadData <= x"0000000000000000";
					when x"8c8" => ReadData <= x"0000000000000000";
					when x"8d0" => ReadData <= x"0000000000000000";
					when x"8d8" => ReadData <= x"0000000000000000";
					when x"8e0" => ReadData <= x"0000000000000000";
					when x"8e8" => ReadData <= x"0000000000000000";
					when x"8f0" => ReadData <= x"0000000000000000";
					when x"8f8" => ReadData <= x"0000000000000000";
					when x"900" => ReadData <= x"0000000000000000";
					when x"908" => ReadData <= x"0000000000000000";
					when x"910" => ReadData <= x"0000000000000000";
					when x"918" => ReadData <= x"0000000000000000";
					when x"920" => ReadData <= x"0000000000000000";
					when x"928" => ReadData <= x"0000000000000000";
					when x"930" => ReadData <= x"0000000000000000";
					when x"938" => ReadData <= x"0000000000000000";
					when x"940" => ReadData <= x"0000000000000000";
					when x"948" => ReadData <= x"0000000000000000";
					when x"950" => ReadData <= x"0000000000000000";
					when x"958" => ReadData <= x"0000000000000000";
					when x"960" => ReadData <= x"0000000000000000";
					when x"968" => ReadData <= x"0000000000000000";
					when x"970" => ReadData <= x"0000000000000000";
					when x"978" => ReadData <= x"0000000000000000";
					when x"980" => ReadData <= x"0000000000000000";
					when x"988" => ReadData <= x"0000000000000000";
					when x"990" => ReadData <= x"0000000000000000";
					when x"998" => ReadData <= x"0000000000000000";
					when x"9a0" => ReadData <= x"0000000000000000";
					when x"9a8" => ReadData <= x"0000000000000000";
					when x"9b0" => ReadData <= x"0000000000000000";
					when x"9b8" => ReadData <= x"0000000000000000";
					when x"9c0" => ReadData <= x"0000000000000000";
					when x"9c8" => ReadData <= x"0000000000000000";
					when x"9d0" => ReadData <= x"0000000000000000";
					when x"9d8" => ReadData <= x"0000000000000000";
					when x"9e0" => ReadData <= x"0000000000000000";
					when x"9e8" => ReadData <= x"0000000000000000";
					when x"9f0" => ReadData <= x"0000000000000000";
					when x"9f8" => ReadData <= x"0000000000000000";
					when x"a00" => ReadData <= x"0000000000000000";
					when x"a08" => ReadData <= x"0000000000000000";
					when x"a10" => ReadData <= x"0000000000000000";
					when x"a18" => ReadData <= x"0000000000000000";
					when x"a20" => ReadData <= x"0000000000000000";
					when x"a28" => ReadData <= x"0000000000000000";
					when x"a30" => ReadData <= x"0000000000000000";
					when x"a38" => ReadData <= x"0000000000000000";
					when x"a40" => ReadData <= x"0000000000000000";
					when x"a48" => ReadData <= x"0000000000000000";
					when x"a50" => ReadData <= x"0000000000000000";
					when x"a58" => ReadData <= x"0000000000000000";
					when x"a60" => ReadData <= x"0000000000000000";
					when x"a68" => ReadData <= x"0000000000000000";
					when x"a70" => ReadData <= x"0000000000000000";
					when x"a78" => ReadData <= x"0000000000000000";
					when x"a80" => ReadData <= x"0000000000000000";
					when x"a88" => ReadData <= x"0000000000000000";
					when x"a90" => ReadData <= x"0000000000000000";
					when x"a98" => ReadData <= x"0000000000000000";
					when x"aa0" => ReadData <= x"0000000000000000";
					when x"aa8" => ReadData <= x"0000000000000000";
					when x"ab0" => ReadData <= x"0000000000000000";
					when x"ab8" => ReadData <= x"0000000000000000";
					when x"ac0" => ReadData <= x"0000000000000000";
					when x"ac8" => ReadData <= x"0000000000000000";
					when x"ad0" => ReadData <= x"0000000000000000";
					when x"ad8" => ReadData <= x"0000000000000000";
					when x"ae0" => ReadData <= x"0000000000000000";
					when x"ae8" => ReadData <= x"0000000000000000";
					when x"af0" => ReadData <= x"0000000000000000";
					when x"af8" => ReadData <= x"0000000000000000";
					when x"b00" => ReadData <= x"0000000000000000";
					when x"b08" => ReadData <= x"0000000000000000";
					when x"b10" => ReadData <= x"0000000000000000";
					when x"b18" => ReadData <= x"0000000000000000";
					when x"b20" => ReadData <= x"0000000000000000";
					when x"b28" => ReadData <= x"0000000000000000";
					when x"b30" => ReadData <= x"0000000000000000";
					when x"b38" => ReadData <= x"0000000000000000";
					when x"b40" => ReadData <= x"0000000000000000";
					when x"b48" => ReadData <= x"0000000000000000";
					when x"b50" => ReadData <= x"0000000000000000";
					when x"b58" => ReadData <= x"0000000000000000";
					when x"b60" => ReadData <= x"0000000000000000";
					when x"b68" => ReadData <= x"0000000000000000";
					when x"b70" => ReadData <= x"0000000000000000";
					when x"b78" => ReadData <= x"0000000000000000";
					when x"b80" => ReadData <= x"0000000000000000";
					when x"b88" => ReadData <= x"0000000000000000";
					when x"b90" => ReadData <= x"0000000000000000";
					when x"b98" => ReadData <= x"0000000000000000";
					when x"ba0" => ReadData <= x"0000000000000000";
					when x"ba8" => ReadData <= x"0000000000000000";
					when x"bb0" => ReadData <= x"0000000000000000";
					when x"bb8" => ReadData <= x"0000000000000000";
					when x"bc0" => ReadData <= x"0000000000000000";
					when x"bc8" => ReadData <= x"0000000000000000";
					when x"bd0" => ReadData <= x"0000000000000000";
					when x"bd8" => ReadData <= x"0000000000000000";
					when x"be0" => ReadData <= x"0000000000000000";
					when x"be8" => ReadData <= x"0000000000000000";
					when x"bf0" => ReadData <= x"0000000000000000";
					when x"bf8" => ReadData <= x"0000000000000000";
					when x"c00" => ReadData <= x"0000000000000000";
					when x"c08" => ReadData <= x"0000000000000000";
					when x"c10" => ReadData <= x"0000000000000000";
					when x"c18" => ReadData <= x"0000000000000000";
					when x"c20" => ReadData <= x"0000000000000000";
					when x"c28" => ReadData <= x"0000000000000000";
					when x"c30" => ReadData <= x"0000000000000000";
					when x"c38" => ReadData <= x"0000000000000000";
					when x"c40" => ReadData <= x"0000000000000000";
					when x"c48" => ReadData <= x"0000000000000000";
					when x"c50" => ReadData <= x"0000000000000000";
					when x"c58" => ReadData <= x"0000000000000000";
					when x"c60" => ReadData <= x"0000000000000000";
					when x"c68" => ReadData <= x"0000000000000000";
					when x"c70" => ReadData <= x"0000000000000000";
					when x"c78" => ReadData <= x"0000000000000000";
					when x"c80" => ReadData <= x"0000000000000000";
					when x"c88" => ReadData <= x"0000000000000000";
					when x"c90" => ReadData <= x"0000000000000000";
					when x"c98" => ReadData <= x"0000000000000000";
					when x"ca0" => ReadData <= x"0000000000000000";
					when x"ca8" => ReadData <= x"0000000000000000";
					when x"cb0" => ReadData <= x"0000000000000000";
					when x"cb8" => ReadData <= x"0000000000000000";
					when x"cc0" => ReadData <= x"0000000000000000";
					when x"cc8" => ReadData <= x"0000000000000000";
					when x"cd0" => ReadData <= x"0000000000000000";
					when x"cd8" => ReadData <= x"0000000000000000";
					when x"ce0" => ReadData <= x"0000000000000000";
					when x"ce8" => ReadData <= x"0000000000000000";
					when x"cf0" => ReadData <= x"0000000000000000";
					when x"cf8" => ReadData <= x"0000000000000000";
					when x"d00" => ReadData <= x"0000000000000000";
					when x"d08" => ReadData <= x"0000000000000000";
					when x"d10" => ReadData <= x"0000000000000000";
					when x"d18" => ReadData <= x"0000000000000000";
					when x"d20" => ReadData <= x"0000000000000000";
					when x"d28" => ReadData <= x"0000000000000000";
					when x"d30" => ReadData <= x"0000000000000000";
					when x"d38" => ReadData <= x"0000000000000000";
					when x"d40" => ReadData <= x"0000000000000000";
					when x"d48" => ReadData <= x"0000000000000000";
					when x"d50" => ReadData <= x"0000000000000000";
					when x"d58" => ReadData <= x"0000000000000000";
					when x"d60" => ReadData <= x"0000000000000000";
					when x"d68" => ReadData <= x"0000000000000000";
					when x"d70" => ReadData <= x"0000000000000000";
					when x"d78" => ReadData <= x"0000000000000000";
					when x"d80" => ReadData <= x"0000000000000000";
					when x"d88" => ReadData <= x"0000000000000000";
					when x"d90" => ReadData <= x"0000000000000000";
					when x"d98" => ReadData <= x"0000000000000000";
					when x"da0" => ReadData <= x"0000000000000000";
					when x"da8" => ReadData <= x"0000000000000000";
					when x"db0" => ReadData <= x"0000000000000000";
					when x"db8" => ReadData <= x"0000000000000000";
					when x"dc0" => ReadData <= x"0000000000000000";
					when x"dc8" => ReadData <= x"0000000000000000";
					when x"dd0" => ReadData <= x"0000000000000000";
					when x"dd8" => ReadData <= x"0000000000000000";
					when x"de0" => ReadData <= x"0000000000000000";
					when x"de8" => ReadData <= x"0000000000000000";
					when x"df0" => ReadData <= x"0000000000000000";
					when x"df8" => ReadData <= x"0000000000000000";
					when x"e00" => ReadData <= x"0000000000000000";
					when x"e08" => ReadData <= x"0000000000000000";
					when x"e10" => ReadData <= x"0000000000000000";
					when x"e18" => ReadData <= x"0000000000000000";
					when x"e20" => ReadData <= x"0000000000000000";
					when x"e28" => ReadData <= x"0000000000000000";
					when x"e30" => ReadData <= x"0000000000000000";
					when x"e38" => ReadData <= x"0000000000000000";
					when x"e40" => ReadData <= x"0000000000000000";
					when x"e48" => ReadData <= x"0000000000000000";
					when x"e50" => ReadData <= x"0000000000000000";
					when x"e58" => ReadData <= x"0000000000000000";
					when x"e60" => ReadData <= x"0000000000000000";
					when x"e68" => ReadData <= x"0000000000000000";
					when x"e70" => ReadData <= x"0000000000000000";
					when x"e78" => ReadData <= x"0000000000000000";
					when x"e80" => ReadData <= x"0000000000000000";
					when x"e88" => ReadData <= x"0000000000000000";
					when x"e90" => ReadData <= x"0000000000000000";
					when x"e98" => ReadData <= x"0000000000000000";
					when x"ea0" => ReadData <= x"0000000000000000";
					when x"ea8" => ReadData <= x"0000000000000000";
					when x"eb0" => ReadData <= x"0000000000000000";
					when x"eb8" => ReadData <= x"0000000000000000";
					when x"ec0" => ReadData <= x"0000000000000000";
					when x"ec8" => ReadData <= x"0000000000000000";
					when x"ed0" => ReadData <= x"0000000000000000";
					when x"ed8" => ReadData <= x"0000000000000000";
					when x"ee0" => ReadData <= x"0000000000000000";
					when x"ee8" => ReadData <= x"0000000000000000";
					when x"ef0" => ReadData <= x"0000000000000000";
					when x"ef8" => ReadData <= x"0000000000000000";
					when x"f00" => ReadData <= x"7f7f7f7f7f7f7f7f";
					when x"f08" => ReadData <= x"8080808080808080";
					when x"f10" => ReadData <= x"0000000000000000";
					when x"f18" => ReadData <= x"0000000000000000";
					when x"f20" => ReadData <= x"0000000000000000";
					when x"f28" => ReadData <= x"0000000000000000";
					when x"f30" => ReadData <= x"0000000000000000";
					when x"f38" => ReadData <= x"0000000000000000";
					when x"f40" => ReadData <= x"0000000000000000";
					when x"f48" => ReadData <= x"0000000000000000";
					when x"f50" => ReadData <= x"0000000000000000";
					when x"f58" => ReadData <= x"0000000000000000";
					when x"f60" => ReadData <= x"0000000000000000";
					when x"f68" => ReadData <= x"0000000000000000";
					when x"f70" => ReadData <= x"0000000000000000";
					when x"f78" => ReadData <= x"0000000000000000";
					when x"f80" => ReadData <= x"0000000000000000";
					when x"f88" => ReadData <= x"0000000000000000";
					when x"f90" => ReadData <= x"0000000000000000";
					when x"f98" => ReadData <= x"0000000000000000";
					when x"fa0" => ReadData <= x"0000000000000000";
					when x"fa8" => ReadData <= x"0000000000000000";
					when x"fb0" => ReadData <= x"0000000000000000";
					when x"fb8" => ReadData <= x"0000000000000000";
					when x"fc0" => ReadData <= x"0000000000000000";
					when x"fc8" => ReadData <= x"0000000000000000";
					when x"fd0" => ReadData <= x"0000000000000000";
					when x"fd8" => ReadData <= x"0000000000000000";
					when x"fe0" => ReadData <= x"0000000000000000";
					when x"fe8" => ReadData <= x"0000000000000000";
					when x"ff0" => ReadData <= x"0000000000000000";
					when others => ReadData <= x"0000000000000000";
                end case;
            end if;
        end if;
    end process;
end rtl;
