-- ***********************************************************************
--              |
-- Title        : Implementation and Optimization of a RISC-V Processor on
--              : a FPGA
--              |
-- Developers   : Hans Jakob Damsgaard, Technical University of Denmark
--              : s163915@student.dtu.dk or hansjakobdamsgaard@gmail.com
--              |
-- Purpose      : This file is a part of a full system implemented as part
--              : of a bachelor's thesis at DTU. The thesis is written in
--              : cooperation with the Institute of Mathematics and
--              : Computer Science.
--              : This entity is a generated ROM containing the bootloader
--              : from the compiler.
--              |
-- Revision     : 1.0   (last updated June 28, 2019)
--              |
-- Available at : https://github.com/hansemandse/RVonFPGA
--              |
-- ***********************************************************************

library IEEE;
use IEEE.std_logic_1164.all;

library work;
use work.includes.all;

entity rom_gen is
    port (
        clk, reset : in std_logic;
        -- Memory interface
        Addr : in std_logic_vector(11 downto 0);
        ReadData : out std_logic_vector(DATA_WIDTH-1 downto 0)
    );
end rom_gen;

architecture rtl of rom_gen is
begin
    process (all)
    begin
        if (rising_edge(clk)) then
            if (reset = '1') then
                ReadData <= (others => '0');
            else
                case (Addr) is
					when x"000" => ReadData <= x"0ac000ef00000513";
					when x"008" => ReadData <= x"0010011b094000ef";
					when x"010" => ReadData <= x"00f1011303011113";
					when x"018" => ReadData <= x"0000119700c11113";
					when x"020" => ReadData <= x"0d0000ef6e418193";
					when x"028" => ReadData <= x"00050067198000ef";
					when x"030" => ReadData <= x"03f51513fff00513";
					when x"038" => ReadData <= x"0005050300350513";
					when x"040" => ReadData <= x"000080670ff57513";
					when x"048" => ReadData <= x"03f51513fff00513";
					when x"050" => ReadData <= x"0005050300250513";
					when x"058" => ReadData <= x"000080670ff57513";
					when x"060" => ReadData <= x"03f51513fff00513";
					when x"068" => ReadData <= x"0007078300350713";
					when x"070" => ReadData <= x"fe078ce30ff7f793";
					when x"078" => ReadData <= x"0005050300150513";
					when x"080" => ReadData <= x"000080670ff57513";
					when x"088" => ReadData <= x"03f79793fff00793";
					when x"090" => ReadData <= x"00a7802300178793";
					when x"098" => ReadData <= x"fff0079300008067";
					when x"0a0" => ReadData <= x"0047879303f79793";
					when x"0a8" => ReadData <= x"0000806700a78023";
					when x"0b0" => ReadData <= x"03f79793fff00793";
					when x"0b8" => ReadData <= x"00a7802300578793";
					when x"0c0" => ReadData <= x"fff0051300008067";
					when x"0c8" => ReadData <= x"0045051303f51513";
					when x"0d0" => ReadData <= x"0ff5751300050503";
					when x"0d8" => ReadData <= x"fff0051300008067";
					when x"0e0" => ReadData <= x"0055051303f51513";
					when x"0e8" => ReadData <= x"0ff5751300050503";
					when x"0f0" => ReadData <= x"000017b700008067";
					when x"0f8" => ReadData <= x"8c87b6838c878713";
					when x"100" => ReadData <= x"fff0079300873703";
					when x"108" => ReadData <= x"03f79793fe010113";
					when x"110" => ReadData <= x"00e13c2300d13823";
					when x"118" => ReadData <= x"01f1051301010613";
					when x"120" => ReadData <= x"0017859300278693";
					when x"128" => ReadData <= x"0ff7771300068703";
					when x"130" => ReadData <= x"00064703fe071ce3";
					when x"138" => ReadData <= x"0016061300e58023";
					when x"140" => ReadData <= x"00578593fea614e3";
					when x"148" => ReadData <= x"0ff6f69300058683";
					when x"150" => ReadData <= x"0007870300478793";
					when x"158" => ReadData <= x"0ff7771300869693";
					when x"160" => ReadData <= x"000186b700d76733";
					when x"168" => ReadData <= x"0007861369f68693";
					when x"170" => ReadData <= x"00c1278300012623";
					when x"178" => ReadData <= x"fef6cae30007879b";
					when x"180" => ReadData <= x"0007879b00c12783";
					when x"188" => ReadData <= x"00e6002300079e63";
					when x"190" => ReadData <= x"00f580230087579b";
					when x"198" => ReadData <= x"030717130017071b";
					when x"1a0" => ReadData <= x"00c1278303075713";
					when x"1a8" => ReadData <= x"00f126230017879b";
					when x"1b0" => ReadData <= x"0007879b00c12783";
					when x"1b8" => ReadData <= x"fb5ff06ffcf6d4e3";
					when x"1c0" => ReadData <= x"f007be03000017b7";
					when x"1c8" => ReadData <= x"f087bf03000017b7";
					when x"1d0" => ReadData <= x"f5010113fff00513";
					when x"1d8" => ReadData <= x"0010029303f51513";
					when x"1e0" => ReadData <= x"0a813423000013b7";
					when x"1e8" => ReadData <= x"09213c230a913023";
					when x"1f0" => ReadData <= x"0941342309313823";
					when x"1f8" => ReadData <= x"07613c2309513023";
					when x"200" => ReadData <= x"0035071307713823";
					when x"208" => ReadData <= x"0791302307813423";
					when x"210" => ReadData <= x"05b1382305a13c23";
					when x"218" => ReadData <= x"0530031300150513";
					when x"220" => ReadData <= x"0390089300900413";
					when x"228" => ReadData <= x"00c0049300010e93";
					when x"230" => ReadData <= x"0020099300100913";
					when x"238" => ReadData <= x"00400a9300300a13";
					when x"240" => ReadData <= x"000f0b93000e0b13";
					when x"248" => ReadData <= x"03c29f938a038393";
					when x"250" => ReadData <= x"0ff7f79300070783";
					when x"258" => ReadData <= x"00050783fe078ce3";
					when x"260" => ReadData <= x"fe6796e30ff7f793";
					when x"268" => ReadData <= x"0ff7f79300070783";
					when x"270" => ReadData <= x"00050c03fe078ce3";
					when x"278" => ReadData <= x"fd0c079b0ffc7c13";
					when x"280" => ReadData <= x"60f466630ff7f793";
					when x"288" => ReadData <= x"0ff7f79300070783";
					when x"290" => ReadData <= x"00050783fe078ce3";
					when x"298" => ReadData <= x"40f8ea630ff7f793";
					when x"2a0" => ReadData <= x"0ff7f693fd07879b";
					when x"2a8" => ReadData <= x"0007078300d10023";
					when x"2b0" => ReadData <= x"fe078ce30ff7f793";
					when x"2b8" => ReadData <= x"0ff7f79300050783";
					when x"2c0" => ReadData <= x"fd07879b3ef8e263";
					when x"2c8" => ReadData <= x"004695930ff7f793";
					when x"2d0" => ReadData <= x"0015959b00b7e5b3";
					when x"2d8" => ReadData <= x"0ff5f59300f100a3";
					when x"2e0" => ReadData <= x"fff5881b08058263";
					when x"2e8" => ReadData <= x"020cdc9302081c93";
					when x"2f0" => ReadData <= x"000e869300110793";
					when x"2f8" => ReadData <= x"000e861301978cb3";
					when x"300" => ReadData <= x"0ff7f79300070783";
					when x"308" => ReadData <= x"00050783fe078ce3";
					when x"310" => ReadData <= x"38f8e2630ff7f793";
					when x"318" => ReadData <= x"0ff7f793fd07879b";
					when x"320" => ReadData <= x"0016061300f60023";
					when x"328" => ReadData <= x"00185c9bfd961ce3";
					when x"330" => ReadData <= x"002e8613001c9c93";
					when x"338" => ReadData <= x"0080006f00cc8cb3";
					when x"340" => ReadData <= x"0006c80300260613";
					when x"348" => ReadData <= x"0048181b0016c783";
					when x"350" => ReadData <= x"0107e7b300f7f793";
					when x"358" => ReadData <= x"0006069300f68023";
					when x"360" => ReadData <= x"0015d593ff9610e3";
					when x"368" => ReadData <= x"fff8069b0005881b";
					when x"370" => ReadData <= x"50c054630006861b";
					when x"378" => ReadData <= x"50f4f463ffe8079b";
					when x"380" => ReadData <= x"000137830036d69b";
					when x"388" => ReadData <= x"00813c8311268863";
					when x"390" => ReadData <= x"0197c7b301c7fd33";
					when x"398" => ReadData <= x"019d0cb301ccfcb3";
					when x"3a0" => ReadData <= x"00fcc7b301e7f7b3";
					when x"3a8" => ReadData <= x"01013c830f368863";
					when x"3b0" => ReadData <= x"00fcc7b301c7fd33";
					when x"3b8" => ReadData <= x"01ac8cb301ccfcb3";
					when x"3c0" => ReadData <= x"00fcc7b301e7f7b3";
					when x"3c8" => ReadData <= x"01813c830d468863";
					when x"3d0" => ReadData <= x"00fcc7b301c7fd33";
					when x"3d8" => ReadData <= x"019d0cb301ccfcb3";
					when x"3e0" => ReadData <= x"00fcc7b301e7f7b3";
					when x"3e8" => ReadData <= x"02013c830b568863";
					when x"3f0" => ReadData <= x"00500d9301c7fd33";
					when x"3f8" => ReadData <= x"01ccfcb30197c7b3";
					when x"400" => ReadData <= x"01e7f7b3019d0cb3";
					when x"408" => ReadData <= x"09b6866300fcc7b3";
					when x"410" => ReadData <= x"01c7fd3302813c83";
					when x"418" => ReadData <= x"0197c7b300600d93";
					when x"420" => ReadData <= x"019d0cb301ccfcb3";
					when x"428" => ReadData <= x"00fcc7b301e7f7b3";
					when x"430" => ReadData <= x"03013c8307b68463";
					when x"438" => ReadData <= x"00700d9301c7fd33";
					when x"440" => ReadData <= x"01ccfcb30197c7b3";
					when x"448" => ReadData <= x"01e7f7b3019d0cb3";
					when x"450" => ReadData <= x"05b6826300fcc7b3";
					when x"458" => ReadData <= x"01c7fd3303813c83";
					when x"460" => ReadData <= x"0197c7b300800d93";
					when x"468" => ReadData <= x"019d0cb301ccfcb3";
					when x"470" => ReadData <= x"00fcc7b301e7f7b3";
					when x"478" => ReadData <= x"0401368303b68063";
					when x"480" => ReadData <= x"00d7c7b30167fcb3";
					when x"488" => ReadData <= x"00dc86b30166f6b3";
					when x"490" => ReadData <= x"00f6c7b30177f7b3";
					when x"498" => ReadData <= x"00f686bb0087d693";
					when x"4a0" => ReadData <= x"00b686bb0107dc93";
					when x"4a8" => ReadData <= x"0187dc93019686bb";
					when x"4b0" => ReadData <= x"0207dc93019686bb";
					when x"4b8" => ReadData <= x"0287dc93019686bb";
					when x"4c0" => ReadData <= x"0307dc93019686bb";
					when x"4c8" => ReadData <= x"0387d793019686bb";
					when x"4d0" => ReadData <= x"ff867c9300f687bb";
					when x"4d8" => ReadData <= x"000c869b0ff7f793";
					when x"4e0" => ReadData <= x"05010c9317960263";
					when x"4e8" => ReadData <= x"fb0ccd0300dc8cb3";
					when x"4f0" => ReadData <= x"00fd07bb00168c9b";
					when x"4f8" => ReadData <= x"14ccd4630ff7f793";
					when x"500" => ReadData <= x"019d0cb305010d13";
					when x"508" => ReadData <= x"00268c9bfb0ccd03";
					when x"510" => ReadData <= x"0ff7f79300fd07bb";
					when x"518" => ReadData <= x"05010d1312ccd663";
					when x"520" => ReadData <= x"fb0ccd03019d0cb3";
					when x"528" => ReadData <= x"00fd07bb00368c9b";
					when x"530" => ReadData <= x"10ccd8630ff7f793";
					when x"538" => ReadData <= x"019d0cb305010d13";
					when x"540" => ReadData <= x"00468c9bfb0ccd03";
					when x"548" => ReadData <= x"0ff7f79300fd07bb";
					when x"550" => ReadData <= x"05010d130eccda63";
					when x"558" => ReadData <= x"fb0ccd03019d0cb3";
					when x"560" => ReadData <= x"00fd07bb00568c9b";
					when x"568" => ReadData <= x"0cccdc630ff7f793";
					when x"570" => ReadData <= x"019d0cb305010d13";
					when x"578" => ReadData <= x"00668c9bfb0ccd03";
					when x"580" => ReadData <= x"0ff7f79300fd07bb";
					when x"588" => ReadData <= x"05010d130accde63";
					when x"590" => ReadData <= x"fb0ccd03019d0cb3";
					when x"598" => ReadData <= x"00fd07bb00768c9b";
					when x"5a0" => ReadData <= x"0accd0630ff7f793";
					when x"5a8" => ReadData <= x"019d0cb305010d13";
					when x"5b0" => ReadData <= x"00868c9bfb0ccd03";
					when x"5b8" => ReadData <= x"0ff7f79300fd07bb";
					when x"5c0" => ReadData <= x"05010d1308ccd263";
					when x"5c8" => ReadData <= x"fb0ccd03019d0cb3";
					when x"5d0" => ReadData <= x"00fd07bb00968c9b";
					when x"5d8" => ReadData <= x"06ccd4630ff7f793";
					when x"5e0" => ReadData <= x"019d0cb305010d13";
					when x"5e8" => ReadData <= x"00a68c9bfb0ccd03";
					when x"5f0" => ReadData <= x"0ff7f79300fd07bb";
					when x"5f8" => ReadData <= x"05010d1304ccd663";
					when x"600" => ReadData <= x"fb0ccd03019d0cb3";
					when x"608" => ReadData <= x"00fd07bb00b68c9b";
					when x"610" => ReadData <= x"02ccd8630ff7f793";
					when x"618" => ReadData <= x"019d0cb305010d13";
					when x"620" => ReadData <= x"00c6869bfb0ccc83";
					when x"628" => ReadData <= x"0ff7f79300fc87bb";
					when x"630" => ReadData <= x"00dd06b300c6da63";
					when x"638" => ReadData <= x"00f687bbfb06c683";
					when x"640" => ReadData <= x"050106930ff7f793";
					when x"648" => ReadData <= x"fb08468301068833";
					when x"650" => ReadData <= x"0ff6f693fff6c693";
					when x"658" => ReadData <= x"fcfc079b24f69063";
					when x"660" => ReadData <= x"008006930ff7f793";
					when x"668" => ReadData <= x"0027979302f6e463";
					when x"670" => ReadData <= x"0007a783007787b3";
					when x"678" => ReadData <= x"0001468300078067";
					when x"680" => ReadData <= x"ffe2879b00114603";
					when x"688" => ReadData <= x"20f6926300c686b3";
					when x"690" => ReadData <= x"bbdff06f0012829b";
					when x"698" => ReadData <= x"0ff7f793fc97879b";
					when x"6a0" => ReadData <= x"fc97879bc81ff06f";
					when x"6a8" => ReadData <= x"c21ff06f0ff7f793";
					when x"6b0" => ReadData <= x"0ff7f693fc97879b";
					when x"6b8" => ReadData <= x"00014503bf1ff06f";
					when x"6c0" => ReadData <= x"0031468300114703";
					when x"6c8" => ReadData <= x"0185151b00214783";
					when x"6d0" => ReadData <= x"00e565330107171b";
					when x"6d8" => ReadData <= x"0087979b00d56533";
					when x"6e0" => ReadData <= x"0005051b00f56533";
					when x"6e8" => ReadData <= x"0a0134830a813403";
					when x"6f0" => ReadData <= x"0901398309813903";
					when x"6f8" => ReadData <= x"08013a8308813a03";
					when x"700" => ReadData <= x"07013b8307813b03";
					when x"708" => ReadData <= x"06013c8306813c03";
					when x"710" => ReadData <= x"05013d8305813d03";
					when x"718" => ReadData <= x"000080670b010113";
					when x"720" => ReadData <= x"0011478300014503";
					when x"728" => ReadData <= x"0105151b00214703";
					when x"730" => ReadData <= x"00f565330087979b";
					when x"738" => ReadData <= x"fadff06f00e56533";
					when x"740" => ReadData <= x"0087d71b00015783";
					when x"748" => ReadData <= x"00e565330087951b";
					when x"750" => ReadData <= x"0305551303051513";
					when x"758" => ReadData <= x"00014803f91ff06f";
					when x"760" => ReadData <= x"00314c0300114683";
					when x"768" => ReadData <= x"0188181b00214783";
					when x"770" => ReadData <= x"00d868330106969b";
					when x"778" => ReadData <= x"0087979b01886833";
					when x"780" => ReadData <= x"0008081b00f86833";
					when x"788" => ReadData <= x"ffa5869bf0cad4e3";
					when x"790" => ReadData <= x"0011079302069693";
					when x"798" => ReadData <= x"00f686b30206d693";
					when x"7a0" => ReadData <= x"000e879341d805b3";
					when x"7a8" => ReadData <= x"0047c80300f58633";
					when x"7b0" => ReadData <= x"0106002301f66633";
					when x"7b8" => ReadData <= x"fed796e300178793";
					when x"7c0" => ReadData <= x"a8dff06f0012829b";
					when x"7c8" => ReadData <= x"0011478300014683";
					when x"7d0" => ReadData <= x"0106969b00214803";
					when x"7d8" => ReadData <= x"00f6e6b30087979b";
					when x"7e0" => ReadData <= x"eaca56e30106e6b3";
					when x"7e8" => ReadData <= x"02059813ffb5859b";
					when x"7f0" => ReadData <= x"0208581300110793";
					when x"7f8" => ReadData <= x"41d685b300f80833";
					when x"800" => ReadData <= x"00f586b3000e8793";
					when x"808" => ReadData <= x"01f6e6b30037c603";
					when x"810" => ReadData <= x"0017879300c68023";
					when x"818" => ReadData <= x"0012829bff0796e3";
					when x"820" => ReadData <= x"00015783a31ff06f";
					when x"828" => ReadData <= x"0087969b0087d81b";
					when x"830" => ReadData <= x"030696930106e6b3";
					when x"838" => ReadData <= x"e4c9dae30306d693";
					when x"840" => ReadData <= x"02059813ffc5859b";
					when x"848" => ReadData <= x"0208581300110793";
					when x"850" => ReadData <= x"41d685b300f80833";
					when x"858" => ReadData <= x"00f586b3000e8793";
					when x"860" => ReadData <= x"01f6e6b30027c603";
					when x"868" => ReadData <= x"0017879300c68023";
					when x"870" => ReadData <= x"0012829bff0796e3";
					when x"878" => ReadData <= x"000587939d9ff06f";
					when x"880" => ReadData <= x"00058793dc5ff06f";
					when x"888" => ReadData <= x"c59ff06f00000693";
					when x"890" => ReadData <= x"e55ff06ffff00513";
					when x"898" => ReadData <= x"e4dff06f00200513";
					when x"8a0" => ReadData <= x"000007c800000824";
					when x"8a8" => ReadData <= x"000006900000075c";
					when x"8b0" => ReadData <= x"000006900000067c";
					when x"8b8" => ReadData <= x"0000072000000740";
					when x"8c0" => ReadData <= x"00000000000006bc";
					when x"8c8" => ReadData <= x"2073692073696854";
					when x"8d0" => ReadData <= x"0021562d43534952";
					when x"8d8" => ReadData <= x"0000000000000000";
					when x"8e0" => ReadData <= x"0000000000000000";
					when x"8e8" => ReadData <= x"0000000000000000";
					when x"8f0" => ReadData <= x"0000000000000000";
					when x"8f8" => ReadData <= x"0000000000000000";
					when x"900" => ReadData <= x"0000000000000000";
					when x"908" => ReadData <= x"0000000000000000";
					when x"910" => ReadData <= x"0000000000000000";
					when x"918" => ReadData <= x"0000000000000000";
					when x"920" => ReadData <= x"0000000000000000";
					when x"928" => ReadData <= x"0000000000000000";
					when x"930" => ReadData <= x"0000000000000000";
					when x"938" => ReadData <= x"0000000000000000";
					when x"940" => ReadData <= x"0000000000000000";
					when x"948" => ReadData <= x"0000000000000000";
					when x"950" => ReadData <= x"0000000000000000";
					when x"958" => ReadData <= x"0000000000000000";
					when x"960" => ReadData <= x"0000000000000000";
					when x"968" => ReadData <= x"0000000000000000";
					when x"970" => ReadData <= x"0000000000000000";
					when x"978" => ReadData <= x"0000000000000000";
					when x"980" => ReadData <= x"0000000000000000";
					when x"988" => ReadData <= x"0000000000000000";
					when x"990" => ReadData <= x"0000000000000000";
					when x"998" => ReadData <= x"0000000000000000";
					when x"9a0" => ReadData <= x"0000000000000000";
					when x"9a8" => ReadData <= x"0000000000000000";
					when x"9b0" => ReadData <= x"0000000000000000";
					when x"9b8" => ReadData <= x"0000000000000000";
					when x"9c0" => ReadData <= x"0000000000000000";
					when x"9c8" => ReadData <= x"0000000000000000";
					when x"9d0" => ReadData <= x"0000000000000000";
					when x"9d8" => ReadData <= x"0000000000000000";
					when x"9e0" => ReadData <= x"0000000000000000";
					when x"9e8" => ReadData <= x"0000000000000000";
					when x"9f0" => ReadData <= x"0000000000000000";
					when x"9f8" => ReadData <= x"0000000000000000";
					when x"a00" => ReadData <= x"0000000000000000";
					when x"a08" => ReadData <= x"0000000000000000";
					when x"a10" => ReadData <= x"0000000000000000";
					when x"a18" => ReadData <= x"0000000000000000";
					when x"a20" => ReadData <= x"0000000000000000";
					when x"a28" => ReadData <= x"0000000000000000";
					when x"a30" => ReadData <= x"0000000000000000";
					when x"a38" => ReadData <= x"0000000000000000";
					when x"a40" => ReadData <= x"0000000000000000";
					when x"a48" => ReadData <= x"0000000000000000";
					when x"a50" => ReadData <= x"0000000000000000";
					when x"a58" => ReadData <= x"0000000000000000";
					when x"a60" => ReadData <= x"0000000000000000";
					when x"a68" => ReadData <= x"0000000000000000";
					when x"a70" => ReadData <= x"0000000000000000";
					when x"a78" => ReadData <= x"0000000000000000";
					when x"a80" => ReadData <= x"0000000000000000";
					when x"a88" => ReadData <= x"0000000000000000";
					when x"a90" => ReadData <= x"0000000000000000";
					when x"a98" => ReadData <= x"0000000000000000";
					when x"aa0" => ReadData <= x"0000000000000000";
					when x"aa8" => ReadData <= x"0000000000000000";
					when x"ab0" => ReadData <= x"0000000000000000";
					when x"ab8" => ReadData <= x"0000000000000000";
					when x"ac0" => ReadData <= x"0000000000000000";
					when x"ac8" => ReadData <= x"0000000000000000";
					when x"ad0" => ReadData <= x"0000000000000000";
					when x"ad8" => ReadData <= x"0000000000000000";
					when x"ae0" => ReadData <= x"0000000000000000";
					when x"ae8" => ReadData <= x"0000000000000000";
					when x"af0" => ReadData <= x"0000000000000000";
					when x"af8" => ReadData <= x"0000000000000000";
					when x"b00" => ReadData <= x"0000000000000000";
					when x"b08" => ReadData <= x"0000000000000000";
					when x"b10" => ReadData <= x"0000000000000000";
					when x"b18" => ReadData <= x"0000000000000000";
					when x"b20" => ReadData <= x"0000000000000000";
					when x"b28" => ReadData <= x"0000000000000000";
					when x"b30" => ReadData <= x"0000000000000000";
					when x"b38" => ReadData <= x"0000000000000000";
					when x"b40" => ReadData <= x"0000000000000000";
					when x"b48" => ReadData <= x"0000000000000000";
					when x"b50" => ReadData <= x"0000000000000000";
					when x"b58" => ReadData <= x"0000000000000000";
					when x"b60" => ReadData <= x"0000000000000000";
					when x"b68" => ReadData <= x"0000000000000000";
					when x"b70" => ReadData <= x"0000000000000000";
					when x"b78" => ReadData <= x"0000000000000000";
					when x"b80" => ReadData <= x"0000000000000000";
					when x"b88" => ReadData <= x"0000000000000000";
					when x"b90" => ReadData <= x"0000000000000000";
					when x"b98" => ReadData <= x"0000000000000000";
					when x"ba0" => ReadData <= x"0000000000000000";
					when x"ba8" => ReadData <= x"0000000000000000";
					when x"bb0" => ReadData <= x"0000000000000000";
					when x"bb8" => ReadData <= x"0000000000000000";
					when x"bc0" => ReadData <= x"0000000000000000";
					when x"bc8" => ReadData <= x"0000000000000000";
					when x"bd0" => ReadData <= x"0000000000000000";
					when x"bd8" => ReadData <= x"0000000000000000";
					when x"be0" => ReadData <= x"0000000000000000";
					when x"be8" => ReadData <= x"0000000000000000";
					when x"bf0" => ReadData <= x"0000000000000000";
					when x"bf8" => ReadData <= x"0000000000000000";
					when x"c00" => ReadData <= x"0000000000000000";
					when x"c08" => ReadData <= x"0000000000000000";
					when x"c10" => ReadData <= x"0000000000000000";
					when x"c18" => ReadData <= x"0000000000000000";
					when x"c20" => ReadData <= x"0000000000000000";
					when x"c28" => ReadData <= x"0000000000000000";
					when x"c30" => ReadData <= x"0000000000000000";
					when x"c38" => ReadData <= x"0000000000000000";
					when x"c40" => ReadData <= x"0000000000000000";
					when x"c48" => ReadData <= x"0000000000000000";
					when x"c50" => ReadData <= x"0000000000000000";
					when x"c58" => ReadData <= x"0000000000000000";
					when x"c60" => ReadData <= x"0000000000000000";
					when x"c68" => ReadData <= x"0000000000000000";
					when x"c70" => ReadData <= x"0000000000000000";
					when x"c78" => ReadData <= x"0000000000000000";
					when x"c80" => ReadData <= x"0000000000000000";
					when x"c88" => ReadData <= x"0000000000000000";
					when x"c90" => ReadData <= x"0000000000000000";
					when x"c98" => ReadData <= x"0000000000000000";
					when x"ca0" => ReadData <= x"0000000000000000";
					when x"ca8" => ReadData <= x"0000000000000000";
					when x"cb0" => ReadData <= x"0000000000000000";
					when x"cb8" => ReadData <= x"0000000000000000";
					when x"cc0" => ReadData <= x"0000000000000000";
					when x"cc8" => ReadData <= x"0000000000000000";
					when x"cd0" => ReadData <= x"0000000000000000";
					when x"cd8" => ReadData <= x"0000000000000000";
					when x"ce0" => ReadData <= x"0000000000000000";
					when x"ce8" => ReadData <= x"0000000000000000";
					when x"cf0" => ReadData <= x"0000000000000000";
					when x"cf8" => ReadData <= x"0000000000000000";
					when x"d00" => ReadData <= x"0000000000000000";
					when x"d08" => ReadData <= x"0000000000000000";
					when x"d10" => ReadData <= x"0000000000000000";
					when x"d18" => ReadData <= x"0000000000000000";
					when x"d20" => ReadData <= x"0000000000000000";
					when x"d28" => ReadData <= x"0000000000000000";
					when x"d30" => ReadData <= x"0000000000000000";
					when x"d38" => ReadData <= x"0000000000000000";
					when x"d40" => ReadData <= x"0000000000000000";
					when x"d48" => ReadData <= x"0000000000000000";
					when x"d50" => ReadData <= x"0000000000000000";
					when x"d58" => ReadData <= x"0000000000000000";
					when x"d60" => ReadData <= x"0000000000000000";
					when x"d68" => ReadData <= x"0000000000000000";
					when x"d70" => ReadData <= x"0000000000000000";
					when x"d78" => ReadData <= x"0000000000000000";
					when x"d80" => ReadData <= x"0000000000000000";
					when x"d88" => ReadData <= x"0000000000000000";
					when x"d90" => ReadData <= x"0000000000000000";
					when x"d98" => ReadData <= x"0000000000000000";
					when x"da0" => ReadData <= x"0000000000000000";
					when x"da8" => ReadData <= x"0000000000000000";
					when x"db0" => ReadData <= x"0000000000000000";
					when x"db8" => ReadData <= x"0000000000000000";
					when x"dc0" => ReadData <= x"0000000000000000";
					when x"dc8" => ReadData <= x"0000000000000000";
					when x"dd0" => ReadData <= x"0000000000000000";
					when x"dd8" => ReadData <= x"0000000000000000";
					when x"de0" => ReadData <= x"0000000000000000";
					when x"de8" => ReadData <= x"0000000000000000";
					when x"df0" => ReadData <= x"0000000000000000";
					when x"df8" => ReadData <= x"0000000000000000";
					when x"e00" => ReadData <= x"0000000000000000";
					when x"e08" => ReadData <= x"0000000000000000";
					when x"e10" => ReadData <= x"0000000000000000";
					when x"e18" => ReadData <= x"0000000000000000";
					when x"e20" => ReadData <= x"0000000000000000";
					when x"e28" => ReadData <= x"0000000000000000";
					when x"e30" => ReadData <= x"0000000000000000";
					when x"e38" => ReadData <= x"0000000000000000";
					when x"e40" => ReadData <= x"0000000000000000";
					when x"e48" => ReadData <= x"0000000000000000";
					when x"e50" => ReadData <= x"0000000000000000";
					when x"e58" => ReadData <= x"0000000000000000";
					when x"e60" => ReadData <= x"0000000000000000";
					when x"e68" => ReadData <= x"0000000000000000";
					when x"e70" => ReadData <= x"0000000000000000";
					when x"e78" => ReadData <= x"0000000000000000";
					when x"e80" => ReadData <= x"0000000000000000";
					when x"e88" => ReadData <= x"0000000000000000";
					when x"e90" => ReadData <= x"0000000000000000";
					when x"e98" => ReadData <= x"0000000000000000";
					when x"ea0" => ReadData <= x"0000000000000000";
					when x"ea8" => ReadData <= x"0000000000000000";
					when x"eb0" => ReadData <= x"0000000000000000";
					when x"eb8" => ReadData <= x"0000000000000000";
					when x"ec0" => ReadData <= x"0000000000000000";
					when x"ec8" => ReadData <= x"0000000000000000";
					when x"ed0" => ReadData <= x"0000000000000000";
					when x"ed8" => ReadData <= x"0000000000000000";
					when x"ee0" => ReadData <= x"0000000000000000";
					when x"ee8" => ReadData <= x"0000000000000000";
					when x"ef0" => ReadData <= x"0000000000000000";
					when x"ef8" => ReadData <= x"0000000000000000";
					when x"f00" => ReadData <= x"7f7f7f7f7f7f7f7f";
					when x"f08" => ReadData <= x"8080808080808080";
					when x"f10" => ReadData <= x"0000000000000000";
					when x"f18" => ReadData <= x"0000000000000000";
					when x"f20" => ReadData <= x"0000000000000000";
					when x"f28" => ReadData <= x"0000000000000000";
					when x"f30" => ReadData <= x"0000000000000000";
					when x"f38" => ReadData <= x"0000000000000000";
					when x"f40" => ReadData <= x"0000000000000000";
					when x"f48" => ReadData <= x"0000000000000000";
					when x"f50" => ReadData <= x"0000000000000000";
					when x"f58" => ReadData <= x"0000000000000000";
					when x"f60" => ReadData <= x"0000000000000000";
					when x"f68" => ReadData <= x"0000000000000000";
					when x"f70" => ReadData <= x"0000000000000000";
					when x"f78" => ReadData <= x"0000000000000000";
					when x"f80" => ReadData <= x"0000000000000000";
					when x"f88" => ReadData <= x"0000000000000000";
					when x"f90" => ReadData <= x"0000000000000000";
					when x"f98" => ReadData <= x"0000000000000000";
					when x"fa0" => ReadData <= x"0000000000000000";
					when x"fa8" => ReadData <= x"0000000000000000";
					when x"fb0" => ReadData <= x"0000000000000000";
					when x"fb8" => ReadData <= x"0000000000000000";
					when x"fc0" => ReadData <= x"0000000000000000";
					when x"fc8" => ReadData <= x"0000000000000000";
					when x"fd0" => ReadData <= x"0000000000000000";
					when x"fd8" => ReadData <= x"0000000000000000";
					when x"fe0" => ReadData <= x"0000000000000000";
					when x"fe8" => ReadData <= x"0000000000000000";
					when x"ff0" => ReadData <= x"0000000000000000";
					when others => ReadData <= x"0000000000000000";
                end case;
            end if;
        end if;
    end process;
end rtl;
